module SimpleReservationStation(
  input         clock,
  input         reset,
  output        io_alloc_ready,
  input         io_alloc_valid,
  input  [1:0]  io_alloc_bits_qType,
  input         io_alloc_bits_opa_valid,
  input  [15:0] io_alloc_bits_opa_start,
  input  [15:0] io_alloc_bits_opa_len,
  input         io_alloc_bits_opb_valid,
  input  [15:0] io_alloc_bits_opb_start,
  input  [15:0] io_alloc_bits_opb_len,
  input         io_alloc_bits_opaIsDst,
  input         io_completed_valid,
  input  [2:0]  io_completed_bits,
  output        io_issue_ld_valid,
  input         io_issue_ld_ready,
  output [1:0]  io_issue_ld_cmd_qType,
  output        io_issue_ld_cmd_opa_valid,
  output [15:0] io_issue_ld_cmd_opa_start,
  output [15:0] io_issue_ld_cmd_opa_len,
  output        io_issue_ld_cmd_opb_valid,
  output [15:0] io_issue_ld_cmd_opb_start,
  output [15:0] io_issue_ld_cmd_opb_len,
  output        io_issue_ld_cmd_opaIsDst,
  output [2:0]  io_issue_ld_robId,
  output        io_issue_ex_valid,
  input         io_issue_ex_ready,
  output [1:0]  io_issue_ex_cmd_qType,
  output        io_issue_ex_cmd_opa_valid,
  output [15:0] io_issue_ex_cmd_opa_start,
  output [15:0] io_issue_ex_cmd_opa_len,
  output        io_issue_ex_cmd_opb_valid,
  output [15:0] io_issue_ex_cmd_opb_start,
  output [15:0] io_issue_ex_cmd_opb_len,
  output        io_issue_ex_cmd_opaIsDst,
  output [2:0]  io_issue_ex_robId,
  output        io_issue_st_valid,
  input         io_issue_st_ready,
  output [1:0]  io_issue_st_cmd_qType,
  output        io_issue_st_cmd_opa_valid,
  output [15:0] io_issue_st_cmd_opa_start,
  output [15:0] io_issue_st_cmd_opa_len,
  output        io_issue_st_cmd_opb_valid,
  output [15:0] io_issue_st_cmd_opb_start,
  output [15:0] io_issue_st_cmd_opb_len,
  output        io_issue_st_cmd_opaIsDst,
  output [2:0]  io_issue_st_robId,
  output        io_busy
);
endmodule
